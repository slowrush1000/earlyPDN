
.SUBCKT INV IN OUT
MN OUT IN VSS VSS N l=10u w=20u
MP OUT IN VDD VDD P l=10u w=30u
R1 IN OUT 1k
.ENDS

.SUBCKT BLOCK IN OUT
XINV1 IN 1 INV
XINV2 2 OUT INV
.ENDS

.SUBCKT TOP IN OUT
XBLOCK1 IN 1 BLOCK
XBLOCK2 2 OUT BLOCK
.ENDS